module Decoder_Pipeline_0(
);
endmodule

module Decoder_Pipeline_1();
endmodule

module Issue_Register_0();
endmodule

module Issue_Register_1();
endmodule

module Branch_Pipeline_Ex();
endmodule

module Memory_Pipeline_Ex();
endmodule

module Branch_Pipeline_Mem();
endmodule

module Memory_Pipeline_Mem();
endmodule

module Branch_Pipeline_WB();
endmodule

module Memory_Pipeline_WB();
endmodule

